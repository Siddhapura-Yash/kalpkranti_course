/* Verilog Implementation of not Gate  */


module m_not (input in,
	    output out);

  assign out = ~in;

endmodule 

